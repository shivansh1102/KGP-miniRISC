`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    15:49:41 10/21/2022 
// Design Name: 
// Module Name:    Diff 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module Diff(input signed[31:0] a, input signed[31:0] b, output reg[31:0] ind);

	wire[31:0] xorAB;
	wire[31:0] onesCompl;
	wire[31:0] compl;
	wire[31:0] ans;

	assign xorAB = a^b;
	assign onesCompl = ~xorAB;

	Adder add3(.a(onesCompl), .b(0), .c_in(1'b1), .sum(compl), .c_out());
	assign ans = xorAB & compl;

	always @(*)
		begin
			case (ans)
				32'b00000000000000000000000000000001: ind = 32'd0;
				32'b00000000000000000000000000000010: ind = 32'd1;
				32'b00000000000000000000000000000100: ind = 32'd2;
				32'b00000000000000000000000000001000: ind = 32'd3;
				32'b00000000000000000000000000010000: ind = 32'd4;
				32'b00000000000000000000000000100000: ind = 32'd5;
				32'b00000000000000000000000001000000: ind = 32'd6;
				32'b00000000000000000000000010000000: ind = 32'd7;
				32'b00000000000000000000000100000000: ind = 32'd8;
				32'b00000000000000000000001000000000: ind = 32'd9;
				32'b00000000000000000000010000000000: ind = 32'd10;
				32'b00000000000000000000100000000000: ind = 32'd11;
				32'b00000000000000000001000000000000: ind = 32'd12;
				32'b00000000000000000010000000000000: ind = 32'd13;
				32'b00000000000000000100000000000000: ind = 32'd14;
				32'b00000000000000001000000000000000: ind = 32'd15;
				32'b00000000000000010000000000000000: ind = 32'd16;
				32'b00000000000000100000000000000000: ind = 32'd17;
				32'b00000000000001000000000000000000: ind = 32'd18;
				32'b00000000000010000000000000000000: ind = 32'd19;
				32'b00000000000100000000000000000000: ind = 32'd20;
				32'b00000000001000000000000000000000: ind = 32'd21;
				32'b00000000010000000000000000000000: ind = 32'd22;
				32'b00000000100000000000000000000000: ind = 32'd23;
				32'b00000001000000000000000000000000: ind = 32'd24;
				32'b00000010000000000000000000000000: ind = 32'd25;
				32'b00000100000000000000000000000000: ind = 32'd26;
				32'b00001000000000000000000000000000: ind = 32'd27;
				32'b00010000000000000000000000000000: ind = 32'd28;
				32'b00100000000000000000000000000000: ind = 32'd29;
				32'b01000000000000000000000000000000: ind = 32'd30;
				32'b10000000000000000000000000000000: ind = 32'd31;
				default: ind = 32'd32;
			endcase
		end

endmodule
